

library ieee;
use ieee.std_logic_1164.all;
use ieee.fixed_pkg.all;
use ieee.math_complex.all;

entity prbs is
end entity prbs;

