

class modem_class;
end modem_class; // UNMATCHED !!

